//====================================================
// Блок регистров FPU процессора PDP2011
//====================================================
module fpuregs (
   input[2:0] raddr,    // адрес чтения
   input[2:0] waddr,    // адрес записи
   input[63:0] d,       // входные данные
   output [63:0] o,     // выходные данные
   input fpmode,        // 0 - 32-битный режим, 1 - 64-битный
   input we,            // строб записи
   input clk            // синхросигнал
);	

// Массив регистров, отдельно старшие и младшие слова
reg[31:0] fpregh[5:0]; // биты 63-32
reg[31:0] fpregl[5:0]; // биты 31-00

//*************************************************
//*  Запись регистров
//*************************************************
always @(posedge clk)  begin
	if (we == 1'b1 & waddr[2:1] != 2'b11)   begin
	   // старшие 32 бита
		fpregh[waddr] <= d[63:32] ; 
		// младшие 32 бита
		if (fpmode == 1'b1) fpregl[waddr] <= d[31:0] ; 
	end  
end 

//*************************************************
//*  Чтение регистров
//*************************************************
assign o = (fpmode == 1'b1)? {fpregh[raddr], fpregl[raddr]} :  // 64-битные данные
			                    {fpregh[raddr], {32{1'b0}}   } ;  // 32-битные данные

endmodule
